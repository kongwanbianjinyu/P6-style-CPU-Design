module testbench;
	// always #5 clk = ~clk;
	
	initial begin
        // $display("value: %d, %d, %d", if_NPC_out[2], if_NPC_out[1], if_NPC_out[0]);
		$finish;
		
	end
	
endmodule